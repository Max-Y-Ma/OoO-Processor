`define EARLY_BRANCH
// `define NORMAL_BRANCH

