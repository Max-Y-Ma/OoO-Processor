`define NUM_TESTS (5000)
