// Top UVM Test Package
`include "frontend_config.svh"

package frontend_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "frontend_sequence.svh"
  `include "frontend_agent.svh"
  `include "frontend_env.svh"
  `include "frontend_test.svh"
endpackage : frontend_pkg
