`define NUM_TESTS (5000)
`define FIFO_WIDTH (32)
`define FIFO_DEPTH (8)